`timescale 1ns / 1ps

module tb;
	
	
	wire count;
	

endmodule